module generators

import strings

const (
	vgen_prelude  = $embed_file('generators/preludes/vgen_v.vfile')
	vgen_postlude = $embed_file('generators/postludes/vgen_v.vfile')
)

/*
** V code Generator
** Why? Because I can.
*/

struct VGenBackend {}

// Generate code for Brainfuck code
fn (cgen VGenBackend) generate_code(options CodeGenInterfaceOptions) ! {
	mut prelude := generators.vgen_prelude.to_string()
	prelude = prelude.replace('mut memory := [255]u8{}', 'mut memory := [${options.memory_size}]u8{}')

	mut output := strings.new_builder(50_000)
	output.write_string('/* Generated by BFCC */\n\n')
	output.write_string(prelude)

	mut indent := 1
	for tok in options.il {
		line := indent_str('\t', indent, match tok.type_token {
			.move_right {
				'ptr += ${tok.value}'
			}
			.move_left {
				'ptr -= ${tok.value}'
			}
			.add {
				'memory[ptr] += ${tok.value}'
			}
			.sub {
				'memory[ptr] -= ${tok.value}'
			}
			.exit {
				'exit(0)'
			}
			.jump_if_zero {
				'for memory[ptr] != 0 {'
			}
			.jump_if_not_zero {
				indent--
				'}'
			}
			.input {
				'memory[ptr] = u8(input_character());'
			}
			.output {
				'print_character(memory[ptr])'
			}
		})
		if tok.type_token == .jump_if_zero {
			indent++
		}
		output.write_string(line)
		output.write_rune(`\n`)
	}

	// Add postlude
	output.write_string(generators.vgen_postlude.to_string())

	// Write to file
	write_code_to_single_file_or_stdout(output.str(), options.output_file, options.print_stdout) or {
		return error('Failed to write code to file')
	}
}
